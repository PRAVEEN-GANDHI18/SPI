`include "/home/ams13/spi/tb/tb1.sv"
