`include "tb1.sv"
